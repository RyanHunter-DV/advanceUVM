module tb;
	initial begin
		$display("hello started");
		#200ns;
		$finish;
	end

endmodule 
