`ifndef uvm_resourceBase__svh
`define uvm_resourceBase__svh


virtual class uvm_resourceBase extends uvm_object; // {

	// scope variable for searching like a hiearachical path
	local string scope;


endclass // }


`endif
