`ifndef regUnit_commandLayer__sv
`define regUnit_commandLayer__sv


class commandLayerClass; // {




endclass // }


`endif
