`ifndef regUnit_regTrans__sv
`define regUnit_regTrans__sv

class regTransClass; // {



endclass // }

`endif
