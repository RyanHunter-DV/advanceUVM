`ifndef smodel_commandBase__sv
`define smodel_commandBase__sv

virtual class commandBaseClass; // {


endclass // }


`endif
