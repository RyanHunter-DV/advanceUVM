`ifndef regUnit_pkg__sv
`define regUnit_pkg__sv

package regUnit; // {

	import smodelBase::*;


endpackage // }


`endif
