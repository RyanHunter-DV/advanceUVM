`ifndef uvm_common__svh
`define uvm_common__svh

`include "common/uvm_types.svh"


`endif
